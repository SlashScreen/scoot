module main 

fn compile_program(input string) ! {
	return error("Todo")
}
