module main


struct Sema {

}
